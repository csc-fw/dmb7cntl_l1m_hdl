`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:07:06 11/19/2015 
// Design Name: 
// Module Name:    trigcon 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module trigcon #(
	parameter TMR = 0
)
(
	input CLK,
	input DRCK,
	input DIN,
	input SEL,
	input FLOAD,
	input FCYC,
	input FCYCM,
	input SHIFT,
	input RST,
	input PLSINJEN,
	input CCBPED,
	output LCTOUT,
	output GTRGOUT
);

wire [1:0] doutl;
wire [13:0] waddr;
wire [12:0] raddr;
//(* ram_style = "block" *)
//reg trig_ram [16383:0];
wire sela;
reg  renb;
reg  cycle;
reg  fcyc_1;
reg  stop;
wire le_fcyc;
wire clr_waddr;
wire clr_raddr;



assign sela = SEL & FLOAD;
assign clr_waddr = !(SHIFT && FLOAD);
assign clr_raddr = (stop || RST);
assign le_fcyc   = FCYC & ~fcyc_1;
assign LCTOUT    = doutl[0];
assign GTRGOUT   = doutl[1];

// Write address counter
cbnce #(
	.Width(14),
	.TMR(TMR)
)
waddr_cnt_i (
	.CLK(DRCK),
	.RST(clr_waddr),
	.CE(1'b1),
	.Q(waddr)
);

// Read address counter
cbnce #(
	.Width(13),
	.TMR(TMR)
)
raddr_cnt_i (
	.CLK(CLK),
	.RST(clr_raddr),
	.CE(renb),
	.Q(raddr)
);

always @(posedge CLK)
begin
	fcyc_1 <= FCYC;
end

always @(posedge CLK or posedge clr_raddr)
begin
	if(clr_raddr)
		cycle <= 1'b0;
	else
		if(CCBPED | le_fcyc)
			cycle <= 1'b1;
end

always @(posedge CLK)
begin
	if(PLSINJEN)
		renb <= cycle | FCYCM;
end

always @(posedge CLK or posedge RST)
begin
	if(RST)
		stop <= 1'b0;
	else
		stop <= raddr[11];
end


//
// Trigger memory
//
//always @(posedge DRCK)
//begin
//	if (sela)
//		if (SHIFT) begin
//			trig_ram[waddr] <= DIN;
//		end
//end
//
//always @(posedge CLK)
//begin
//	if (RST)
//		doutl <= 2'b00;
//	if (renb)
//		begin
//			doutl[0] <= trig_ram[{raddr, 1'b0}];
//			doutl[1] <= trig_ram[{raddr, 1'b1}];
//		end
//end



   // RAMB16_S1_S2: Virtex-II/II-Pro, Spartan-3/3E 16k/8k x 1/2 Dual-Port RAM
   // Xilinx HDL Language Template, version 10.1.3

   RAMB16_S1_S2 #(
      .INIT_A(1'b0),   // Value of output RAM registers on Port A at startup
      .INIT_B(2'b00),  // Value of output RAM registers on Port B at startup
      .SRVAL_A(1'b0),  // Port A output value upon SSR assertion
      .SRVAL_B(2'b00), // Port B output value upon SSR assertion
      .WRITE_MODE_A("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .WRITE_MODE_B("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE
      .SIM_COLLISION_CHECK("ALL"),  // "NONE", "WARNING_ONLY", "GENERATE_X_ONLY", "ALL" 

      // The following INIT_xx declarations specify the initial contents of the RAM
      // Port A Address 0 to 4095, Port B Address 0 to 2047
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Port A Address 4096 to 8191, Port B Address 2048 to 4095
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Port A Address 8192 to 12287, Port B Address 4095 to 6143
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Port A Address 12288 to 16383, Port B Address 6144 to 8091 
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000)
   ) RAMB16_S1_S2_inst (
      .DOA(),         // Port A 1-bit Data Output
      .DOB(doutl),    // Port B 2-bit Data Output
      .ADDRA(waddr),  // Port A 14-bit Address Input
      .ADDRB(raddr),  // Port B 13-bit Address Input
      .CLKA(DRCK),    // Port A Clock
      .CLKB(CLK),     // Port B Clock
      .DIA(DIN),      // Port A 1-bit Data Input
      .DIB(2'b0),     // Port B 2-bit Data Input
      .ENA(sela),     // Port A RAM Enable Input
      .ENB(renb),     // Port B RAM Enable Input
      .SSRA(RST),     // Port A Synchronous Set/Reset Input
      .SSRB(RST),     // Port B Synchronous Set/Reset Input
      .WEA(SHIFT),    // Port A Write Enable Input
      .WEB(1'b0)      // Port B Write Enable Input
   );

endmodule
